magic
tech tsmc
timestamp 1755744555
<< nwell >>
rect -15 0 28 25
rect 38 -1 95 25
rect 133 -1 190 25
rect 37 -92 94 -66
rect 132 -92 189 -66
<< ntransistor >>
rect 5 -39 9 -29
rect 56 -38 60 -29
rect 73 -38 77 -29
rect 151 -38 155 -29
rect 168 -38 172 -29
rect 55 -129 59 -120
rect 72 -129 76 -120
rect 150 -129 154 -120
rect 167 -129 171 -120
<< ptransistor >>
rect 5 8 9 17
rect 56 8 60 17
rect 73 8 77 17
rect 151 8 155 17
rect 168 8 172 17
rect 55 -83 59 -74
rect 72 -83 76 -74
rect 150 -83 154 -74
rect 167 -83 171 -74
<< ndiffusion >>
rect -7 -30 5 -29
rect -7 -38 -5 -30
rect 3 -38 5 -30
rect -7 -39 5 -38
rect 9 -30 20 -29
rect 9 -38 11 -30
rect 19 -38 20 -30
rect 54 -37 56 -29
rect 46 -38 56 -37
rect 60 -38 73 -29
rect 77 -37 79 -29
rect 87 -37 88 -29
rect 77 -38 88 -37
rect 149 -37 151 -29
rect 141 -38 151 -37
rect 155 -38 168 -29
rect 172 -37 174 -29
rect 182 -37 183 -29
rect 172 -38 183 -37
rect 9 -39 20 -38
rect 53 -128 55 -120
rect 45 -129 55 -128
rect 59 -129 72 -120
rect 76 -128 78 -120
rect 86 -128 87 -120
rect 76 -129 87 -128
rect 148 -128 150 -120
rect 140 -129 150 -128
rect 154 -129 167 -120
rect 171 -128 173 -120
rect 181 -128 182 -120
rect 171 -129 182 -128
<< pdiffusion >>
rect -7 9 -5 17
rect 3 9 5 17
rect -7 8 5 9
rect 9 9 11 17
rect 19 9 20 17
rect 9 8 20 9
rect 54 9 56 17
rect 46 8 56 9
rect 60 9 62 17
rect 70 9 73 17
rect 60 8 73 9
rect 77 9 79 17
rect 77 8 87 9
rect 149 9 151 17
rect 141 8 151 9
rect 155 9 157 17
rect 165 9 168 17
rect 155 8 168 9
rect 172 9 174 17
rect 172 8 182 9
rect 53 -82 55 -74
rect 45 -83 55 -82
rect 59 -82 61 -74
rect 69 -82 72 -74
rect 59 -83 72 -82
rect 76 -82 78 -74
rect 76 -83 86 -82
rect 148 -82 150 -74
rect 140 -83 150 -82
rect 154 -82 156 -74
rect 164 -82 167 -74
rect 154 -83 167 -82
rect 171 -82 173 -74
rect 171 -83 181 -82
<< ndcontact >>
rect -5 -38 3 -30
rect 11 -38 19 -30
rect 46 -37 54 -29
rect 79 -37 87 -29
rect 141 -37 149 -29
rect 174 -37 182 -29
rect 45 -128 53 -120
rect 78 -128 86 -120
rect 140 -128 148 -120
rect 173 -128 181 -120
<< pdcontact >>
rect -5 9 3 17
rect 11 9 19 17
rect 46 9 54 17
rect 62 9 70 17
rect 79 9 87 17
rect 141 9 149 17
rect 157 9 165 17
rect 174 9 182 17
rect 45 -82 53 -74
rect 61 -82 69 -74
rect 78 -82 86 -74
rect 140 -82 148 -74
rect 156 -82 164 -74
rect 173 -82 181 -74
<< psubstratepcontact >>
rect 11 -52 19 -44
rect 46 -52 54 -44
rect 141 -52 149 -44
rect 45 -143 53 -135
rect 140 -143 148 -135
<< nsubstratencontact >>
rect 11 25 19 33
rect 58 25 67 33
rect 153 25 162 33
rect 57 -66 66 -58
rect 152 -66 161 -58
<< polysilicon >>
rect 5 17 9 21
rect 56 17 60 21
rect 73 17 77 21
rect 151 17 155 21
rect 168 17 172 21
rect 5 -7 9 8
rect 56 -7 60 8
rect -29 -15 -9 -10
rect -29 -108 -23 -15
rect 5 -13 60 -7
rect 5 -29 9 -13
rect 56 -29 60 -13
rect 73 -2 77 8
rect 73 -10 74 -2
rect 73 -29 77 -10
rect 151 -15 155 8
rect 90 -22 155 -15
rect 151 -29 155 -22
rect 168 -4 172 8
rect 168 -7 205 -4
rect 168 -29 172 -7
rect 185 -22 195 -15
rect 5 -43 9 -39
rect 56 -42 60 -38
rect 73 -42 77 -38
rect 151 -42 155 -38
rect 168 -42 172 -38
rect 55 -74 59 -70
rect 72 -74 76 -70
rect 150 -74 154 -70
rect 167 -74 171 -70
rect 55 -108 59 -83
rect -29 -113 59 -108
rect 55 -120 59 -113
rect 72 -93 76 -83
rect 72 -101 73 -93
rect 72 -120 76 -101
rect 150 -106 154 -83
rect 89 -113 154 -106
rect 150 -120 154 -113
rect 167 -95 171 -83
rect 192 -95 195 -22
rect 167 -99 195 -95
rect 167 -120 171 -99
rect 200 -106 205 -7
rect 184 -113 205 -106
rect 55 -133 59 -129
rect 72 -133 76 -129
rect 150 -133 154 -129
rect 167 -133 171 -129
<< polycontact >>
rect -9 -17 -1 -9
rect 74 -10 82 -2
rect 82 -23 90 -15
rect 177 -23 185 -15
rect 73 -101 81 -93
rect 81 -114 89 -106
rect 176 -114 184 -106
<< metal1 >>
rect 19 25 58 33
rect 67 25 153 33
rect 162 25 213 33
rect 11 17 19 25
rect 46 17 54 25
rect 79 17 87 25
rect 141 17 149 25
rect 174 17 182 25
rect -5 -9 3 9
rect -1 -17 3 -9
rect -5 -30 3 -17
rect 62 -15 70 9
rect 82 -9 107 -4
rect 62 -22 82 -15
rect 79 -23 82 -22
rect 79 -29 87 -23
rect 11 -44 19 -38
rect 100 -27 107 -9
rect 157 -15 165 9
rect 157 -22 177 -15
rect 46 -44 54 -37
rect 174 -23 177 -22
rect 174 -29 182 -23
rect 19 -52 46 -45
rect 141 -44 149 -37
rect 54 -52 141 -45
rect 149 -52 179 -44
rect 11 -135 19 -52
rect 207 -58 213 25
rect 45 -66 57 -58
rect 66 -66 152 -58
rect 161 -66 213 -58
rect 45 -74 53 -66
rect 78 -74 86 -66
rect 61 -106 69 -82
rect 140 -74 148 -66
rect 173 -74 181 -66
rect 100 -95 107 -83
rect 81 -99 107 -95
rect 156 -106 164 -82
rect 61 -113 81 -106
rect 78 -114 81 -113
rect 156 -113 176 -106
rect 173 -114 176 -113
rect 78 -120 86 -114
rect 173 -120 181 -114
rect 45 -135 53 -128
rect 140 -135 148 -128
rect 11 -143 45 -135
rect 53 -143 140 -135
rect 148 -143 151 -135
<< m2contact >>
rect 100 -41 107 -27
rect 100 -83 107 -72
<< metal2 >>
rect 100 -72 107 -41
<< labels >>
rlabel polysilicon 76 -12 76 -12 1 clk
rlabel metal1 110 30 110 30 5 vdd
rlabel polysilicon 46 -9 46 -9 1 D
rlabel polysilicon 188 -17 188 -17 1 q
rlabel metal1 101 -138 101 -138 1 Gnd
rlabel polysilicon 194 -110 194 -110 1 q_bar
<< end >>
